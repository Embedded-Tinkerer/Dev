module registers (clk, CE, D, Q);


endmodule